module alu(input [15:0]A, B, input [3:0] shift_amt, opcode,
		output [15:0] S, output N, Z, V);



endmodule